module Final_Project();

		NES_driver inst();


endmodule