module Final_Project();

		NES_driver inst();
		PS2_Controller inst2();

endmodule